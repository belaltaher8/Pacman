module sum_1la(a, b, cin, s);

	input a, b, cin;
	output s;

	xor xor0(s, a, b, cin);


endmodule